//这是QamCarrier.v文件的程序清单
module QamCarrier (
	rst,clk,din,
	di,dq,df); 
	
	input		rst;   //复位信号，高电平有效
	input		clk;   //时钟信号，数据速率/采样速率/FPGA系统时钟/8 MHz
	input	 signed [7:0]	din;    //输入的16QAM已调数据
	output signed [26:0]	di;     //解调后的基带信号(同相支路)
	output signed [26:0]	dq;     //解调后的基带信号(正交支路)
	output signed [26:0]	df;     //环路滤波器输出数据
	
	//首先对输入数据通过寄存器输入
   /*	
	reg signed [7:0] din1,dint;
	always @(posedge clk or posedge rst)
	   if (rst)
		   begin
			   din1 <= 8'd0;
				dint <= 8'd0;
			end
		else
	      begin
			   din1 <= din;
				dint <= din1;
			end
	*/
	reg signed [7:0] dint;
	always @(posedge clk)
	   dint <= din;
	
	//实例化NCO核所需的接口信号
	wire reset_n,out_valid,clken;
	wire [30:0] carrier;
	wire signed [9:0] sin,cos ;
	wire signed [30:0] frequency_df;
	wire signed [26:0] Loopout;
	assign reset_n = !rst;
	assign clken = 1'b1;
	assign carrier=31'd536870912;//2MHz  df=0Hz
	//assign carrier=31'd537005130;//2.0005MHz  df=500Hz
	//assign carrier=31'd537139347;//2.001MHz   df=1KHz
	assign frequency_df={{4{Loopout[26]}},Loopout};//根据NCO核接口，扩展为30位
	
	//实例化NCO核
   //Quartus提供的NCO核输出数据最小位宽为10比特，根据环路设计需求，只取高8比特参与后续运算	
	nco	u0 (
		.phi_inc_i (carrier),
		.clk (clk),
		.reset_n (reset_n),
		.clken (clken),
		.freq_mod_i (frequency_df),
		.fsin_o (sin),
		.fcos_o (cos),
		.out_valid (out_valid));
	
   //实例化NCO同相支路乘法运算器核
	wire signed [15:0] zi;	
   mult8_8 u1 (
	   .clock (clk),
		.dataa (sin[9:2]),
		.datab (dint),
		.result (zi));
		
   //实例化NCO正交支路乘法运算器核	
	wire signed [15:0] zq;	
   mult8_8 u2 (
	   .clock (clk),
		.dataa (cos[9:2]),
		.datab (dint),
		.result (zq));
		

   //实例化鉴相器同相支路低通滤波器核
	wire ast_sink_valid,ast_source_ready;
	wire [1:0] ast_sink_error;
	assign ast_sink_valid=1'b1;
	assign ast_source_ready=1'b1;
	assign ast_sink_error=2'd0;
	wire sink_readyi,source_validi;
	wire [1:0] source_errori;
	wire signed [26:0] yi;	
   fir_lpf u3(
		.clk (clk),
		.reset_n (reset_n),
		.ast_sink_data (zi[14:0]),
		.ast_sink_valid (ast_sink_valid),
		.ast_source_ready (ast_source_ready),
		.ast_sink_error (ast_sink_error),
		.ast_source_data (yi),
		.ast_sink_ready (sink_readyi),
		.ast_source_valid (source_validi),
		.ast_source_error (source_errori));


   //实例化鉴相器正交支路低通滤波器核
	wire sink_readyq,source_validq;
	wire [1:0] source_errorq;
	wire signed [26:0] yq;	
   fir_lpf u4(
		.clk (clk),
		.reset_n (reset_n),
		.ast_sink_data (zq[14:0]),
		.ast_sink_valid (ast_sink_valid),
		.ast_source_ready (ast_source_ready),
		.ast_sink_error (ast_sink_error),
		.ast_source_data (yq),
		.ast_sink_ready (sink_readyq),
		.ast_source_valid (source_validq),
		.ast_source_error (source_errorq));
		
		
	//实例化鉴相器模块
	wire signed [26:0] pd;
	PolarDetect u6 (
	   .rst (rst),
		.clk (clk),
		.yi (yi),
		.yq (yq),
		.pd (pd));
			
	//实例化环路滤波器模块	
   LoopFilter u5(
	   .rst (rst),
		.clk (clk),
		.pd  (pd),
		.frequency_df(Loopout));
		

   //对时钟分频，产生位同步模块时钟信号clk_half
	reg clk_half;
	reg signed [15:0] dig,dqg;

	always @(posedge clk or posedge rst)
	   if (rst)
		   begin
		      clk_half <= 1'b0;
				dig <= 16'd0;
				dqg <= 16'd0;
			end
		else
		   begin
		      clk_half <= !clk_half;
				//对基带解调数据实现2倍抽取，送入位同步模块
				if (!clk_half)
				   begin
					   dig <= yi[26:11];
						dqg <= yq[26:11];
					end
			end
			
	wire signed [17:0] yig,yqg;	
	wire signed [15:0] u,e,w;		
	//实例化位同步模块	
   FpgaGardner u7(
	   .rst (rst),
		.clk (clk_half),
		.di  (dig),
		.dq  (dqg),
		.yi  (yig),
		.yq  (yqg),		
		.u(u),
		.e(e),
		.w(w),
		.sync(bitsync));		
		
	
   //匹配滤波后的数据为同相、正交基带信号输出
	assign df = Loopout;
	assign di = {yig,9'd0};
	assign dq = {yqg,9'd0};

	
endmodule
